/*
module cpu_fsm

endmodule
*/

module top_cpu

    
    //Instantiate Instruction memory

    //Instantiate Micro-instruction memory interface

    //Instantiate Register File 


endmodule