module mcontrol #(
    
) (
    sys_clk,
    
);
    
endmodule